configuration io_ctrl_rtl_cfg of io_ctrl is
  for rtl      -- architecture rtl is used for entity io_ctrl
  end for;
end io_ctrl_rtl_cfg;
