-------------------------------------------------------------------------------
-- VGA CONTROLLER PROJECT
-------------------------------------------------------------------------------
-- Author: Konstantin Haferl
--
-- Filename: mem_ctrl_3_.vhd
--
-- Date of Creation: 2023 11 15
--
-- Version: 1.0
--
-- Design Unit: Memory Controller 3 (Testbench)
--
-- Description: The Memory Controller 3 is part of the VGA controller project.
-- The Memory Controller 3 generates addresses for a ROM where a 100x100x12bit
-- image is stored.
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_mem_ctrl_3 is
end tb_mem_ctrl_3;

