-------------------------------------------------------------------------------
--                                                                      
--                        adder_8bit task
--  
-------------------------------------------------------------------------------
--                                                                      
-- ENTITY:         tb_adder_8bit
--
-- FILENAME:       tb_adder_8bit_.vhd
-- 
-- ARCHITECTURE:   sim
-- 
-- ENGINEER:       Konstantin Haferl
--
-- DATE:           20.3.2023
--
-- VERSION:        1.0
--
-------------------------------------------------------------------------------
--                                                                      
-- DESCRIPTION:    This is the entity declaration of the adder_8bit testbench
--                 for the adder_8bit task.
--
-------------------------------------------------------------------------------
--
-- REFERENCES:     (none)
--
-------------------------------------------------------------------------------
--                                                                      
-- PACKAGES:       std_logic_1164 (IEEE library)
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_adder_8bit is
end tb_adder_8bit;

