-------------------------------------------------------------------------------
-- VGA CONTROLLER PROJECT
-------------------------------------------------------------------------------
-- Author: Konstantin Haferl
--
-- Filename: mem_ctrl_2_.vhd
--
-- Date of Creation: 2023 11 13
--
-- Version: 1.0
--
-- Design Unit: Memory Controller 2 (Testbench)
--
-- Description: The Memory Controller 2 is part of the VGA controller project.
-- The Memory Controller 2 generates addresses for a ROM where a 100x100x12bit
-- image is stored.
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_mem_ctrl_2 is
end tb_mem_ctrl_2;

