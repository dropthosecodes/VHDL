-------------------------------------------------------------------------------
--                                                                      
--                        D_FF task
--  
-------------------------------------------------------------------------------
--                                                                      
-- ENTITY:         D_FF
--
-- FILENAME:       D_FF_rtl_cfg.vhd
-- 
-- ARCHITECTURE:   rtl
-- 
-- ENGINEER:       Konstantin Haferl
--
-- DATE:           13.03.2023
--
-- VERSION:        1.0
--
-------------------------------------------------------------------------------
--                                                                      
-- DESCRIPTION:    This is the configuration for the entity D_FF and the
--                 architecture rtl.
--
-------------------------------------------------------------------------------
--
-- REFERENCES:     (none)
--
-------------------------------------------------------------------------------
--                                                                      
-- PACKAGES:       std_logic_1164 (IEEE library)
--
-------------------------------------------------------------------------------

configuration D_FF_rtl_cfg of D_FF is
  for rtl        -- architecture rtl is used for entity D_FF
  end for;
end D_FF_rtl_cfg;
