library IEEE;
use IEEE.std_logic_1164.all;

entity tb_gate_model is
end tb_gate_model;

