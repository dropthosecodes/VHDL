library IEEE;
use IEEE.std_logic_1164.all;

entity tb_led_fsm is
end tb_led_fsm;

