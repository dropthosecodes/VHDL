-------------------------------------------------------------------------------
-- VGA CONTROLLER PROJECT
-------------------------------------------------------------------------------
-- Author: Konstantin Haferl
--
-- Filename: tb_src_mux_.vhd
--
-- Date of Creation: 2023 10 10
--
-- Version: 1.0
--
-- Design Unit: Source Multiplexer (Testbench)
--
-- Description: The Source Multiplexer is part of the VGA controller project.
-- It routes the RGB signals to the VGA Control Unit according to the
-- position of the switches on the Basys3 devboard .
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_src_mux is
end tb_src_mux;

