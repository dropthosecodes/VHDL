configuration mem_ctrl_2_rtl_cfg of mem_ctrl_2 is
  for rtl      -- architecture rtl is used for entity mem_ctrl_2
  end for;
end mem_ctrl_2_rtl_cfg;
