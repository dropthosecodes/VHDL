-------------------------------------------------------------------------------
--                                                                      
--                        adder_8bit task
--  
-------------------------------------------------------------------------------
--                                                                      
-- ENTITY:         adder_8bit
--
-- FILENAME:       adder_8bit_rtl_cfg.vhd
-- 
-- ARCHITECTURE:   rtl
-- 
-- ENGINEER:       Konstantin Haferl
--
-- DATE:           20.03.2023
--
-- VERSION:        1.0
--
-------------------------------------------------------------------------------
--                                                                      
-- DESCRIPTION:    This is the configuration for the entity adder_8bit and the
--                 architecture rtl.
--
-------------------------------------------------------------------------------
--
-- REFERENCES:     (none)
--
-------------------------------------------------------------------------------
--                                                                      
-- PACKAGES:       std_logic_1164 (IEEE library)
--
-------------------------------------------------------------------------------

configuration adder_8bit_rtl_cfg of adder_8bit is
  for rtl        -- architecture rtl is used for entity adder_8bit
  end for;
end adder_8bit_rtl_cfg;
