-- MC8051 IP Core Demo Design, Top-level Configuration
-- FPGA device/board: Xilinx Artix-7 on Digilent Basys3 board
-- Author: Peter Roessler
-- Date: 2017-02-08

configuration fpga_top_rtl_cfg of fpga_top is
    for rtl
    end for;
end fpga_top_rtl_cfg;
