configuration alu_rtl_cfg of alu is
  for rtl      -- architecture rtl is used for entity alu
  end for;
end alu_rtl_cfg;