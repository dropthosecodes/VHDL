configuration pattern_gen_1_rtl_cfg of pattern_gen_1 is
  for rtl      -- architecture rtl is used for entity pattern_gen_1
  end for;
end pattern_gen_1_rtl_cfg;
