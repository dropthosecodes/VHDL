-- MC8051 IP Core Demo Design, Entity for Top-level Testbench 
-- Author: Peter Roessler
-- Date: 2017-02-08

library ieee;
use ieee.std_logic_1164.all;

use std.textio.all;

entity tb_mc8051 is
end;
