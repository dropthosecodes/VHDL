-------------------------------------------------------------------------------
--                                                                      
--                        decoder_3bit task
--  
-------------------------------------------------------------------------------
--                                                                      
-- ENTITY:         decoder_3bit
--
-- FILENAME:       decoder_3bit_rtl_cfg.vhd
-- 
-- ARCHITECTURE:   rtl
-- 
-- ENGINEER:       Konstantin Haferl
--
-- DATE:           27.2.2023
--
-- VERSION:        1.0
--
-------------------------------------------------------------------------------
--                                                                      
-- DESCRIPTION:    This is the configuration for the entity decoder_3bit and the
--                 architecture rtl.
--
-------------------------------------------------------------------------------
--
-- REFERENCES:     (none)
--
-------------------------------------------------------------------------------
--                                                                      
-- PACKAGES:       std_logic_1164 (IEEE library)
--
-------------------------------------------------------------------------------

configuration decoder_3bit_rtl_cfg of decoder_3bit is
  for rtl        -- architecture rtl is used for entity decoder_3bit
  end for;
end decoder_3bit_rtl_cfg;
