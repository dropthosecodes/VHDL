configuration vga_ctrl_rtl_cfg of vga_ctrl is
  for rtl      -- architecture rtl is used for entity vga_ctrl
  end for;
end vga_ctrl_rtl_cfg;
