-- MC8051 IP Core Demo Design, Configuration for Top-level Testbench 
-- Author: Peter Roessler
-- Date: 2017-02-08

configuration tb_mc8051_sim_cfg of tb_mc8051 is
  for sim
  end for;
end tb_mc8051_sim_cfg;
