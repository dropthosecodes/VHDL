configuration mem_ctrl_3_rtl_cfg of mem_ctrl_3 is
  for rtl      -- architecture rtl is used for entity mem_ctrl_3
  end for;
end mem_ctrl_3_rtl_cfg;
