-------------------------------------------------------------------------------
--                                                                      
--                        decoder_3bit task
--  
-------------------------------------------------------------------------------
--                                                                      
-- ENTITY:         tb_decoder_3bit
--
-- FILENAME:       tb_decoder_3bit_.vhd
-- 
-- ARCHITECTURE:   sim
-- 
-- ENGINEER:       Konstantin Haferl
--
-- DATE:           27.2.2023
--
-- VERSION:        1.0
--
-------------------------------------------------------------------------------
--                                                                      
-- DESCRIPTION:    This is the entity declaration of the decoder_3bit testbench
--                 for the decoder_3bit task.
--
-------------------------------------------------------------------------------
--
-- REFERENCES:     (none)
--
-------------------------------------------------------------------------------
--                                                                      
-- PACKAGES:       std_logic_1164 (IEEE library)
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_decoder_3bit is
end tb_decoder_3bit;

