-------------------------------------------------------------------------------
--                                                                      
--                        simplegate task
--  
-------------------------------------------------------------------------------
--                                                                      
-- ENTITY:         tb_xorgate
--
-- FILENAME:       tb_xorgate_.vhd
-- 
-- ARCHITECTURE:   sim
-- 
-- ENGINEER:       Konstantin Haferl
--
-- DATE:           20.2.2023
--
-- VERSION:        1.0
--
-------------------------------------------------------------------------------
--                                                                      
-- DESCRIPTION:    This is the entity declaration of the xorgate testbench
--                 for the simplegate task.
--
-------------------------------------------------------------------------------
--
-- REFERENCES:     (none)
--
-------------------------------------------------------------------------------
--                                                                      
-- PACKAGES:       std_logic_1164 (IEEE library)
--
-------------------------------------------------------------------------------
--                                                                      
-- CHANGES:        Version 1.0 - KH - 20.2.2023
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_xorgate is
end tb_xorgate;

