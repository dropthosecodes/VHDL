configuration train_fsm_rtl_cfg of train_fsm is
  for rtl      -- architecture rtl is used for entity train_fsm
  end for;
end train_fsm_rtl_cfg;
