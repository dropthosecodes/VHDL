configuration prescaler_rtl_cfg of prescaler is
  for rtl      -- architecture rtl is used for entity prescaler
  end for;
end prescaler_rtl_cfg;
