configuration calc_top_struc_cfg of calc_top is
  for struc     -- architecture rtl is used for entity calc_top
  end for;
end calc_top_struc_cfg;
