-------------------------------------------------------------------------------
-- VGA CONTROLLER PROJECT
-------------------------------------------------------------------------------
-- Author: Konstantin Haferl
--
-- Filename: tb_pattern_gen_1_.vhd
--
-- Date of Creation: 2023 09 19
--
-- Version: 1.0
--
-- Design Unit: Pattern Generator 1 (Testbench)
--
-- Description: The Pattern Generator 1 is part of the VGA controller project.
-- It generates a pattern of Red-Green-Blue-Black columns on the 640x480 screen.
-- The columns are 40 pixels wide, therefore a total of 16 columns are generated.
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_pattern_gen_1 is
end tb_pattern_gen_1;

