-------------------------------------------------------------------------------
-- VGA CONTROLLER PROJECT
-------------------------------------------------------------------------------
-- Author: Konstantin Haferl
--
-- Filename: tb_io_logic_.vhd
--
-- Date of Creation: 2023 09 19
--
-- Version: 1.0
--
-- Design Unit: IO Logic Unit (Testbench)
--
-- Description: The IO Logic Unit is part of the VGA controller project
-- It handles the debouncing of the push buttons as well as the three switches SW0, SW1 and SW2.
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_io_logic is
end tb_io_logic;

