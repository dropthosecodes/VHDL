configuration pattern_gen_2_rtl_cfg of pattern_gen_2 is
  for rtl      -- architecture rtl is used for entity pattern_gen_2
  end for;
end pattern_gen_2_rtl_cfg;
