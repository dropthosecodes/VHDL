configuration src_mux_rtl_cfg of src_mux is
  for rtl      -- architecture rtl is used for entity src_mux
  end for;
end src_mux_rtl_cfg;
