-------------------------------------------------------------------------------
-- VGA CONTROLLER PROJECT
-------------------------------------------------------------------------------
-- Author: Konstantin Haferl
--
-- Filename: tb_vga_ctrl_.vhd
--
-- Date of Creation: 2023 09 18
--
-- Version: 1.0
--
-- Design Unit: VGA Control Unit (Testbench)
--
-- Description: The VGA Control unit is part of the VGA controller project
-- It drives the VGA signals and generates the horizontal any vertical sync
-- counters for the memory controllers and pattern generators
--
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_vga_ctrl is
end tb_vga_ctrl;

