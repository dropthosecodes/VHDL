configuration io_logic_rtl_cfg of io_logic is
  for rtl      -- architecture rtl is used for entity io_logic
  end for;
end io_logic_rtl_cfg;
