configuration shift_reg_rtl_cfg of shift_reg is
  for rtl        -- architecture rtl is used for entity shift_reg
  end for;
end shift_reg_rtl_cfg;
