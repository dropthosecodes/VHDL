configuration mem_ctrl_1_rtl_cfg of mem_ctrl_1 is
  for rtl      -- architecture rtl is used for entity mem_ctrl_1
  end for;
end mem_ctrl_1_rtl_cfg;
