library IEEE;
use IEEE.std_logic_1164.all;

entity tb_train_fsm is
end tb_train_fsm;

