-------------------------------------------------------------------------------
--                                                                      
--                        vectorgates task
--  
-------------------------------------------------------------------------------
--                                                                      
-- ENTITY:         tb_vectorgates
--
-- FILENAME:       tb_vectorgates_.vhd
-- 
-- ARCHITECTURE:   sim
-- 
-- ENGINEER:       Konstantin Haferl
--
-- DATE:           27.2.2023
--
-- VERSION:        1.0
--
-------------------------------------------------------------------------------
--                                                                      
-- DESCRIPTION:    This is the entity declaration of the vectorgates testbench
--                 for the vectorgates task.
--
-------------------------------------------------------------------------------
--
-- REFERENCES:     (none)
--
-------------------------------------------------------------------------------
--                                                                      
-- PACKAGES:       std_logic_1164 (IEEE library)
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_vectorgates is
end tb_vectorgates;

