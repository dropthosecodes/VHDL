library IEEE;
use IEEE.std_logic_1164.all;

entity tb_shift_reg is
end tb_shift_reg;

