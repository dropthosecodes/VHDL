-------------------------------------------------------------------------------
-- VGA CONTROLLER PROJECT
-------------------------------------------------------------------------------
-- Author: Konstantin Haferl
--
-- Filename: tb_top_.vhd
--
-- Date of Creation: 2023 11 06
--
-- Version: 1.0
--
-- Design Unit: Top-Level Design of the VGA Controller (Testbench)
--
-- Description: This is the top-level design of the VGA Controller project.
-- It interconnects all sub-units and interfaces to the circuitry of the
-- Digilent Basys3 FPGA board.
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_top is
end tb_top;

