-------------------------------------------------------------------------------
--                                                                      
--                        vectorgates task
--  
-------------------------------------------------------------------------------
--                                                                      
-- ENTITY:         vectorgates
--
-- FILENAME:       vectorgates_rtl_cfg.vhd
-- 
-- ARCHITECTURE:   rtl
-- 
-- ENGINEER:       Konstantin Haferl
--
-- DATE:           27.2.2023
--
-- VERSION:        1.0
--
-------------------------------------------------------------------------------
--                                                                      
-- DESCRIPTION:    This is the configuration for the entity vectorgates and the
--                 architecture rtl.
--
-------------------------------------------------------------------------------
--
-- REFERENCES:     (none)
--
-------------------------------------------------------------------------------
--                                                                      
-- PACKAGES:       std_logic_1164 (IEEE library)
--
-------------------------------------------------------------------------------

configuration vectorgates_rtl_cfg of vectorgates is
  for rtl        -- architecture rtl is used for entity vectorgates
  end for;
end vectorgates_rtl_cfg;
