-------------------------------------------------------------------------------
--                                                                      
--                        JK_FF task
--  
-------------------------------------------------------------------------------
--                                                                      
-- ENTITY:         tb_JK_FF
--
-- FILENAME:       tb_JK_FF_.vhd
-- 
-- ARCHITECTURE:   sim
-- 
-- ENGINEER:       Konstantin Haferl
--
-- DATE:           13.3.2023
--
-- VERSION:        1.0
--
-------------------------------------------------------------------------------
--                                                                      
-- DESCRIPTION:    This is the entity declaration of the JK_FF testbench
--                 for the JK_FF task.
--
-------------------------------------------------------------------------------
--
-- REFERENCES:     (none)
--
-------------------------------------------------------------------------------
--                                                                      
-- PACKAGES:       std_logic_1164 (IEEE library)
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_JK_FF is
end tb_JK_FF;

