-------------------------------------------------------------------------------
--                                                                      
--                        JK_FF task
--  
-------------------------------------------------------------------------------
--                                                                      
-- ENTITY:         JK_FF
--
-- FILENAME:       JK_FF_rtl_cfg.vhd
-- 
-- ARCHITECTURE:   rtl
-- 
-- ENGINEER:       Konstantin Haferl
--
-- DATE:           13.03.2023
--
-- VERSION:        1.0
--
-------------------------------------------------------------------------------
--                                                                      
-- DESCRIPTION:    This is the configuration for the entity JK_FF and the
--                 architecture rtl.
--
-------------------------------------------------------------------------------
--
-- REFERENCES:     (none)
--
-------------------------------------------------------------------------------
--                                                                      
-- PACKAGES:       std_logic_1164 (IEEE library)
--
-------------------------------------------------------------------------------

configuration JK_FF_rtl_cfg of JK_FF is
  for rtl        -- architecture rtl is used for entity JK_FF
  end for;
end JK_FF_rtl_cfg;
