configuration led_fsm_rtl_cfg of led_fsm is
  for rtl        -- architecture rtl is used for entity led_fsm
  end for;
end led_fsm_rtl_cfg;
