configuration vga_controller_top_struc_cfg of vga_controller_top is
  for struc     -- architecture rtl is used for entity vga_controller_top
  end for;
end vga_controller_top_struc_cfg;
